module Reg_Div(init,in_ld,ld,Sub_res,shift_bit,clk);
